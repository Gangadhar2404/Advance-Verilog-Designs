module eqz(in,out);
  input in;
  output out;
  assign out=(in==0);
  endmodule